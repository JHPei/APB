`define D_WIDTH 32
`define MEM_DEPTH 10
`define SLAVE_SUPPD 2
